`ifndef HEEPSILON_CLOCK_CONFIG_SVH
`define HEEPSILON_CLOCK_CONFIG_SVH
`define HEEPSILON_CPU_CLK_HZ 100000000
`define HEEPSILON_CPU_CLK_KHZ 100000
`define HEEPSILON_CGRA_CLK_HZ 100000000
`define HEEPSILON_CGRA_CLK_KHZ 100000
`endif
